/*#########################################################################
#File Name:     ls42_tb.sv
#Description:   SN74LS42 - 4-Line BCD to 10-Line Decimal Decoder test bench.
#                            
#Date:          
#Programmer:    Jonathon McEllin, S00150412
#Version:       Rev. 1.00
#
#Notes:         
##########################################################################*/

`timescale 1ps / 1ps
module ls42_tb; 
/*-------------------------- Inputs and Outputs --------------------------*/
	reg    _A, _B, _C, _D;
 	wire   _0, _1, _2, _3, _4, _5, _6, _7, _8, _9;
	
	
/*--------------------- Instantiate Device Under Test --------------------*/
	ls42 DUT( 
		._A(_A),
		._B(_B),
		._C(_C),
		._D(_D),
		._0(_0),
		._1(_1),
		._2(_2),
		._3(_3),
		._4(_4),
		._5(_5),
		._6(_6),
		._7(_7),
		._8(_8),
		._9(_9)
	);	
		
/*--------------------------------- Test ---------------------------------*/
	initial begin
		_D= 1'b0; _C = 1'b0; _B= 1'b0; _A = 1'b0;
		#0 $display("_A = %b, _B = %b, _C = %b, _D = %b", _A, _B, _C, _D);
		#0 $display("_0 = %b, _1 = %b, _2 = %b, _3 = %b, _4 = %b, _5 = %b, _6 = %b, _7 = %b, _8 = %b, _9 = %b", _0, _1, _2, _3, _4, _5, _6, _7, _8, _9);

		#10 _D= 1'b0; _C = 1'b0; _B= 1'b0; _A = 1'b1;
		#0 $display("_D = %b, _C = %b, _B = %b, _A = %b", _D, _C, _B, _A);
		#0 $display("_0 = %b, _1 = %b, _2 = %b, _3 = %b, _4 = %b, _5 = %b, _6 = %b, _7 = %b, _8 = %b, _9 = %b", _0, _1, _2, _3, _4, _5, _6, _7, _8, _9);

		#10 _D= 1'b0; _C = 1'b0; _B= 1'b1; _A = 1'b0;
		#0 $display("_A = %b, _B = %b, _C = %b, _D = %b", _A, _B, _C, _D);
		#0 $display("_0 = %b, _1 = %b, _2 = %b, _3 = %b, _4 = %b, _5 = %b, _6 = %b, _7 = %b, _8 = %b, _9 = %b", _0, _1, _2, _3, _4, _5, _6, _7, _8, _9);

		#10 _D= 1'b0; _C = 1'b0; _B= 1'b1; _A = 1'b1;
		#0 $display("_D = %b, _C = %b, _B = %b, _A = %b", _D, _C, _B, _A);
		#0 $display("_0 = %b, _1 = %b, _2 = %b, _3 = %b, _4 = %b, _5 = %b, _6 = %b, _7 = %b, _8 = %b, _9 = %b", _0, _1, _2, _3, _4, _5, _6, _7, _8, _9);

		#10 _D= 1'b0; _C = 1'b1; _B= 1'b0; _A = 1'b0;
		#0 $display("_A = %b, _B = %b, _C = %b, _D = %b", _A, _B, _C, _D);
		#0 $display("_0 = %b, _1 = %b, _2 = %b, _3 = %b, _4 = %b, _5 = %b, _6 = %b, _7 = %b, _8 = %b, _9 = %b", _0, _1, _2, _3, _4, _5, _6, _7, _8, _9);

		#10 _D= 1'b0; _C = 1'b1; _B= 1'b0; _A = 1'b1;
		#0 $display("_D = %b, _C = %b, _B = %b, _A = %b", _D, _C, _B, _A);
		#0 $display("_0 = %b, _1 = %b, _2 = %b, _3 = %b, _4 = %b, _5 = %b, _6 = %b, _7 = %b, _8 = %b, _9 = %b", _0, _1, _2, _3, _4, _5, _6, _7, _8, _9);

		#10 _D= 1'b0; _C = 1'b1; _B= 1'b1; _A = 1'b0;
		#0 $display("_A = %b, _B = %b, _C = %b, _D = %b", _A, _B, _C, _D);
		#0 $display("_0 = %b, _1 = %b, _2 = %b, _3 = %b, _4 = %b, _5 = %b, _6 = %b, _7 = %b, _8 = %b, _9 = %b", _0, _1, _2, _3, _4, _5, _6, _7, _8, _9);

		#10 _D= 1'b0; _C = 1'b1; _B= 1'b1; _A = 1'b1;
		#0 $display("_D = %b, _C = %b, _B = %b, _A = %b", _D, _C, _B, _A);
		#0 $display("_0 = %b, _1 = %b, _2 = %b, _3 = %b, _4 = %b, _5 = %b, _6 = %b, _7 = %b, _8 = %b, _9 = %b", _0, _1, _2, _3, _4, _5, _6, _7, _8, _9);

		#10 _D= 1'b1; _C = 1'b0; _B= 1'b0; _A = 1'b0;
		#0 $display("_A = %b, _B = %b, _C = %b, _D = %b", _A, _B, _C, _D);
		#0 $display("_0 = %b, _1 = %b, _2 = %b, _3 = %b, _4 = %b, _5 = %b, _6 = %b, _7 = %b, _8 = %b, _9 = %b", _0, _1, _2, _3, _4, _5, _6, _7, _8, _9);

		#10 _D= 1'b1; _C = 1'b0; _B= 1'b0; _A = 1'b1;
		#0 $display("_D = %b, _C = %b, _B = %b, _A = %b", _D, _C, _B, _A);
		#0 $display("_0 = %b, _1 = %b, _2 = %b, _3 = %b, _4 = %b, _5 = %b, _6 = %b, _7 = %b, _8 = %b, _9 = %b", _0, _1, _2, _3, _4, _5, _6, _7, _8, _9);

		#10 _D= 1'b1; _C = 1'b0; _B= 1'b1; _A = 1'b0;
		#0 $display("_A = %b, _B = %b, _C = %b, _D = %b", _A, _B, _C, _D);
		#0 $display("_0 = %b, _1 = %b, _2 = %b, _3 = %b, _4 = %b, _5 = %b, _6 = %b, _7 = %b, _8 = %b, _9 = %b", _0, _1, _2, _3, _4, _5, _6, _7, _8, _9);

		#10 _D= 1'b1; _C = 1'b0; _B= 1'b1; _A = 1'b1;
		#0 $display("_D = %b, _C = %b, _B = %b, _A = %b", _D, _C, _B, _A);
		#0 $display("_0 = %b, _1 = %b, _2 = %b, _3 = %b, _4 = %b, _5 = %b, _6 = %b, _7 = %b, _8 = %b, _9 = %b", _0, _1, _2, _3, _4, _5, _6, _7, _8, _9);

		#10 _D= 1'b1; _C = 1'b1; _B= 1'b0; _A = 1'b0;
		#0 $display("_A = %b, _B = %b, _C = %b, _D = %b", _A, _B, _C, _D);
		#0 $display("_0 = %b, _1 = %b, _2 = %b, _3 = %b, _4 = %b, _5 = %b, _6 = %b, _7 = %b, _8 = %b, _9 = %b", _0, _1, _2, _3, _4, _5, _6, _7, _8, _9);

		#10 _D= 1'b1; _C = 1'b1; _B= 1'b0; _A = 1'b1;
		#0 $display("_D = %b, _C = %b, _B = %b, _A = %b", _D, _C, _B, _A);
		#0 $display("_0 = %b, _1 = %b, _2 = %b, _3 = %b, _4 = %b, _5 = %b, _6 = %b, _7 = %b, _8 = %b, _9 = %b", _0, _1, _2, _3, _4, _5, _6, _7, _8, _9);

		#10 _D= 1'b1; _C = 1'b1; _B= 1'b1; _A = 1'b0;
		#0 $display("_A = %b, _B = %b, _C = %b, _D = %b", _A, _B, _C, _D);
		#0 $display("_0 = %b, _1 = %b, _2 = %b, _3 = %b, _4 = %b, _5 = %b, _6 = %b, _7 = %b, _8 = %b, _9 = %b", _0, _1, _2, _3, _4, _5, _6, _7, _8, _9);

		#10 _D= 1'b1; _C = 1'b1; _B= 1'b1; _A = 1'b1;
		#0 $display("_D = %b, _C = %b, _B = %b, _A = %b", _D, _C, _B, _A);
		#0 $display("_0 = %b, _1 = %b, _2 = %b, _3 = %b, _4 = %b, _5 = %b, _6 = %b, _7 = %b, _8 = %b, _9 = %b", _0, _1, _2, _3, _4, _5, _6, _7, _8, _9);

		#10 $stop;
	end
	
endmodule