/*#########################################################################
#File Name:     video_playfield.sv
#Description:   Representation of Playfield (Dynamic RAM A) schematic 
#               diagram contained in Kangaroo Schematic Package Supplement 
#				Sheet 11A.
#				 			          
#Date:          
#Programmer:    Jonathon McEllin, S00150412
#Version:       Rev. 1.00
#
#Notes:         
##########################################################################*/

module video_playfield(
	/*-------------------------------------------------------------- /
	/ --------------------- Inputs and Outputs --------------------- /
	/ --------------------------------------------------------------*/
	
	/* -> Playfield */
	input wire SEL_I_II_AL_A,
	input wire AV6_TICK_AL,
	input wire ENA,
	input wire SFT_AL,

	input wire ACAS0_AL,
	input wire ACAS1_AL,
	input wire ARAS0_AL,
	input wire ARAS1_AL,
	input wire AWE0_AL,
	input wire AWE1_AL,

	input wire XXA6,
	input wire XXA5,
	input wire XXA4,
	input wire XXA3,
	input wire XXA2,
	input wire XXA1,
	input wire XXA0,

	input wire DXR3,
	input wire DXR2,
	input wire DXR1,
	input wire DXR0,
	input wire DXG3,
	input wire DXG2,
	input wire DXG1,
	input wire DXG0,
	input wire DXB3,
	input wire DXB2,
	input wire DXB1,
	input wire DXB0,
	input wire DXZ3,
	input wire DXZ2,
	input wire DXZ1,
	input wire DXZ0,

	input wire KOS1,
	input wire ARHF_AL,
	input wire AGHF_AL,
	input wire ABHF_AL,
	input wire BY_AL,
	input wire PRIA_AL,

	output wire AVR,
	output wire AVG,
	output wire AVB,
	output wire AY_AL,
	output wire LD_SFT_AL,
	

	/* -> External Shared Logic */
	/* IC117 - LS04 */
	input wire IC117_10_TO_IC107_1_AND_IC108_1_AND_IC109_1_AND_IC110_1,

	/* IC139 - LS00 */
	input wire IC139_8_TO_IC107_15_AND_IC108_15_AND_IC109_15_AND_IC110_15,
	input wire IC139_11_TO_IC137_2_AND_IC137_3_AND_IC137_11
);


	/*-------------------------------------------------------------- /
	/ --------------------- Nets and Registers --------------------- /
	/-------------------------------------------------------------- */

	/* -> Playfield */
	wire AR, AG, AB, AZ;
	wire IC55_14_TO_IC110_3_AND_IC110_14, IC56_14_TO_IC110_6_AND_IC110_11, IC57_14_TO_IC110_5_AND_IC110_10, IC58_14_TO_IC110_2_AND_IC110_13, IC66_14_TO_IC109_3_AND_IC109_14, IC67_14_TO_IC109_6_AND_IC109_11, IC68_14_TO_IC109_5_AND_IC109_10, IC69_14_TO_IC109_2_AND_IC109_13, IC79_14_TO_IC108_3_AND_IC108_14, IC80_14_TO_IC108_6_AND_IC108_11, IC81_14_TO_IC108_5_AND_IC108_10, IC82_14_TO_IC108_2_AND_IC108_13, IC93_14_TO_IC107_3_AND_IC107_14, IC94_14_TO_IC107_6_AND_IC107_11, IC95_14_TO_IC107_5_AND_IC107_10, IC96_14_TO_IC107_2_AND_IC107_13, IC107_4_TO_IC121_5, IC107_7_TO_IC121_4, IC107_9_TO_IC121_3, IC107_12_TO_IC121_2, IC108_4_TO_IC122_5, IC108_7_TO_IC122_4, IC108_9_TO_IC122_3, IC108_12_TO_IC122_2, IC109_4_TO_IC123_5, IC109_7_TO_IC123_4, IC109_9_TO_IC123_3, IC109_12_TO_IC123_2, IC110_4_TO_IC124_5, IC110_7_TO_IC124_4, IC110_9_TO_IC124_3, IC110_12_TO_IC124_2, IC138_8_TO_IC136_2_AND_IC136_5_AND_IC136_10, IC136_3_TO_IC137_13, IC136_6_TO_IC137_5, IC136_8_TO_IC137_9, IC138_3_TO_IC138_4, IC138_11_TO_IC138_5;


	/*-------------------------------------------------------------- /
	/ --------------------- Module Instantiation ------------------- /
	/ --------------------------------------------------------------*/

	/* -> Playfield */
	/* IC55 - 4116 */
	_4116 IC55(.RAS(ARAS1_AL), .CAS(ACAS1_AL), .WE(AWE1_AL), .A0(XXA0), .A1(XXA1), .A2(XXA2), .A3(XXA3), .A4(XXA4), .A5(XXA5), .A6(XXA6), .D(DXB3), .Q(IC55_14_TO_IC110_3_AND_IC110_14));

	/* IC56 - 4116 */
	_4116 IC56(.RAS(ARAS1_AL), .CAS(ACAS1_AL), .WE(AWE1_AL), .A0(XXA0), .A1(XXA1), .A2(XXA2), .A3(XXA3), .A4(XXA4), .A5(XXA5), .A6(XXA6), .D(DXB2), .Q(IC56_14_TO_IC110_6_AND_IC110_11));

	/* IC57 - 4116 */
	_4116 IC57(.RAS(ARAS1_AL), .CAS(ACAS1_AL), .WE(AWE1_AL), .A0(XXA0), .A1(XXA1), .A2(XXA2), .A3(XXA3), .A4(XXA4), .A5(XXA5), .A6(XXA6), .D(DXB1), .Q(IC57_14_TO_IC110_5_AND_IC110_10));

	/* IC58 - 4116 */
	_4116 IC58(.RAS(ARAS1_AL), .CAS(ACAS1_AL), .WE(AWE1_AL), .A0(XXA0), .A1(XXA1), .A2(XXA2), .A3(XXA3), .A4(XXA4), .A5(XXA5), .A6(XXA6), .D(DXB0), .Q(IC58_14_TO_IC110_2_AND_IC110_13));

	/* IC66 - 4116 */
	_4116 IC66(.RAS(ARAS1_AL), .CAS(ACAS1_AL), .WE(AWE1_AL), .A0(XXA0), .A1(XXA1), .A2(XXA2), .A3(XXA3), .A4(XXA4), .A5(XXA5), .A6(XXA6), .D(DXG3), .Q(IC66_14_TO_IC109_3_AND_IC109_14));

	/* IC67 - 4116 */
	_4116 IC67(.RAS(ARAS1_AL), .CAS(ACAS1_AL), .WE(AWE1_AL), .A0(XXA0), .A1(XXA1), .A2(XXA2), .A3(XXA3), .A4(XXA4), .A5(XXA5), .A6(XXA6), .D(DXG2), .Q(IC67_14_TO_IC109_6_AND_IC109_11));

	/* IC68 - 4116 */
	_4116 IC68(.RAS(ARAS1_AL), .CAS(ACAS1_AL), .WE(AWE1_AL), .A0(XXA0), .A1(XXA1), .A2(XXA2), .A3(XXA3), .A4(XXA4), .A5(XXA5), .A6(XXA6), .D(DXG1), .Q(IC68_14_TO_IC109_5_AND_IC109_10));

	/* IC69 - 4116 */
	_4116 IC69(.RAS(ARAS1_AL), .CAS(ACAS1_AL), .WE(AWE1_AL), .A0(XXA0), .A1(XXA1), .A2(XXA2), .A3(XXA3), .A4(XXA4), .A5(XXA5), .A6(XXA6), .D(DXG0), .Q(IC69_14_TO_IC109_2_AND_IC109_13));

	/* IC79 - 4116 */
	_4116 IC79(.RAS(ARAS0_AL), .CAS(ACAS0_AL), .WE(AWE0_AL), .A0(XXA0), .A1(XXA1), .A2(XXA2), .A3(XXA3), .A4(XXA4), .A5(XXA5), .A6(XXA6), .D(DXR3), .Q(IC79_14_TO_IC108_3_AND_IC108_14));

	/* IC80 - 4116 */
	_4116 IC80(.RAS(ARAS0_AL), .CAS(ACAS0_AL), .WE(AWE0_AL), .A0(XXA0), .A1(XXA1), .A2(XXA2), .A3(XXA3), .A4(XXA4), .A5(XXA5), .A6(XXA6), .D(DXR2), .Q(IC80_14_TO_IC108_6_AND_IC108_11));

	/* IC81 - 4116 */
	_4116 IC81(.RAS(ARAS0_AL), .CAS(ACAS0_AL), .WE(AWE0_AL), .A0(XXA0), .A1(XXA1), .A2(XXA2), .A3(XXA3), .A4(XXA4), .A5(XXA5), .A6(XXA6), .D(DXR1), .Q(IC81_14_TO_IC108_5_AND_IC108_10));

	/* IC82 - 4116 */
	_4116 IC82(.RAS(ARAS0_AL), .CAS(ACAS0_AL), .WE(AWE0_AL), .A0(XXA0), .A1(XXA1), .A2(XXA2), .A3(XXA3), .A4(XXA4), .A5(XXA5), .A6(XXA6), .D(DXR0), .Q(IC82_14_TO_IC108_2_AND_IC108_13));

	/* IC93 - 4116 */
	_4116 IC93(.RAS(ARAS0_AL), .CAS(ACAS0_AL), .WE(AWE0_AL), .A0(XXA0), .A1(XXA1), .A2(XXA2), .A3(XXA3), .A4(XXA4), .A5(XXA5), .A6(XXA6), .D(DXZ3), .Q(IC93_14_TO_IC107_3_AND_IC107_14));

	/* IC94 - 4116 */
	_4116 IC94(.RAS(ARAS0_AL), .CAS(ACAS0_AL), .WE(AWE0_AL), .A0(XXA0), .A1(XXA1), .A2(XXA2), .A3(XXA3), .A4(XXA4), .A5(XXA5), .A6(XXA6), .D(DXZ2), .Q(IC94_14_TO_IC107_6_AND_IC107_11));

	/* IC95 - 4116 */
	_4116 IC95(.RAS(ARAS0_AL), .CAS(ACAS0_AL), .WE(AWE0_AL), .A0(XXA0), .A1(XXA1), .A2(XXA2), .A3(XXA3), .A4(XXA4), .A5(XXA5), .A6(XXA6), .D(DXZ1), .Q(IC95_14_TO_IC107_5_AND_IC107_10));

	/* IC96 - 4116 */
	_4116 IC96(.RAS(ARAS0_AL), .CAS(ACAS0_AL), .WE(AWE0_AL), .A0(XXA0), .A1(XXA1), .A2(XXA2), .A3(XXA3), .A4(XXA4), .A5(XXA5), .A6(XXA6), .D(DXZ0), .Q(IC96_14_TO_IC107_2_AND_IC107_13));

	/* IC107 - LS157 */
	ls157 IC107(._AB(IC117_10_TO_IC107_1_AND_IC108_1_AND_IC109_1_AND_IC110_1), ._G(IC139_8_TO_IC107_15_AND_IC108_15_AND_IC109_15_AND_IC110_15), ._1A(IC96_14_TO_IC107_2_AND_IC107_13), ._1B(IC93_14_TO_IC107_3_AND_IC107_14), ._1Y(IC107_4_TO_IC121_5), ._2A(IC95_14_TO_IC107_5_AND_IC107_10), ._2B(IC94_14_TO_IC107_6_AND_IC107_11), ._2Y(IC107_7_TO_IC121_4), ._3A(IC94_14_TO_IC107_6_AND_IC107_11), ._3B(IC95_14_TO_IC107_5_AND_IC107_10), ._3Y(IC107_9_TO_IC121_3), ._4A(IC93_14_TO_IC107_3_AND_IC107_14), ._4B(IC96_14_TO_IC107_2_AND_IC107_13), ._4Y(IC107_12_TO_IC121_2));

	/* IC108 - LS157 */
	ls157 IC108(._AB(IC117_10_TO_IC107_1_AND_IC108_1_AND_IC109_1_AND_IC110_1), ._G(IC139_8_TO_IC107_15_AND_IC108_15_AND_IC109_15_AND_IC110_15), ._1A(IC82_14_TO_IC108_2_AND_IC108_13), ._1B(IC79_14_TO_IC108_3_AND_IC108_14), ._1Y(IC108_4_TO_IC122_5), ._2A(IC81_14_TO_IC108_5_AND_IC108_10), ._2B(IC80_14_TO_IC108_6_AND_IC108_11), ._2Y(IC108_7_TO_IC122_4), ._3A(IC80_14_TO_IC108_6_AND_IC108_11), ._3B(IC81_14_TO_IC108_5_AND_IC108_10), ._3Y(IC108_9_TO_IC122_3), ._4A(IC79_14_TO_IC108_3_AND_IC108_14), ._4B(IC82_14_TO_IC108_2_AND_IC108_13), ._4Y(IC108_12_TO_IC122_2));

	/* IC109 - LS157 */
	ls157 IC109(._AB(IC117_10_TO_IC107_1_AND_IC108_1_AND_IC109_1_AND_IC110_1), ._G(IC139_8_TO_IC107_15_AND_IC108_15_AND_IC109_15_AND_IC110_15), ._1A(IC69_14_TO_IC109_2_AND_IC109_13), ._1B(IC66_14_TO_IC109_3_AND_IC109_14), ._1Y(IC109_4_TO_IC123_5), ._2A(IC68_14_TO_IC109_5_AND_IC109_10), ._2B(IC67_14_TO_IC109_6_AND_IC109_11), ._2Y(IC109_7_TO_IC123_4), ._3A(IC67_14_TO_IC109_6_AND_IC109_11), ._3B(IC68_14_TO_IC109_5_AND_IC109_10), ._3Y(IC109_9_TO_IC123_3), ._4A(IC66_14_TO_IC109_3_AND_IC109_14), ._4B(IC69_14_TO_IC109_2_AND_IC109_13), ._4Y(IC109_12_TO_IC123_2));

	/* IC110 - LS157 */
	ls157 IC110(._AB(IC117_10_TO_IC107_1_AND_IC108_1_AND_IC109_1_AND_IC110_1), ._G(IC139_8_TO_IC107_15_AND_IC108_15_AND_IC109_15_AND_IC110_15), ._1A(IC58_14_TO_IC110_2_AND_IC110_13), ._1B(IC55_14_TO_IC110_3_AND_IC110_14), ._1Y(IC110_4_TO_IC124_5), ._2A(IC57_14_TO_IC110_5_AND_IC110_10), ._2B(IC56_14_TO_IC110_6_AND_IC110_11), ._2Y(IC110_7_TO_IC124_4), ._3A(IC56_14_TO_IC110_6_AND_IC110_11), ._3B(IC57_14_TO_IC110_5_AND_IC110_10), ._3Y(IC110_9_TO_IC124_3), ._4A(IC55_14_TO_IC110_3_AND_IC110_14), ._4B(IC58_14_TO_IC110_2_AND_IC110_13), ._4Y(IC110_12_TO_IC124_2));

	/* IC121 - LS95 */
	ls95 IC121(._CLK1(SFT_AL), ._CLK2(SFT_AL), ._SER(), ._MODE(LD_SFT_AL), ._A(IC107_12_TO_IC121_2), ._B(IC107_9_TO_IC121_3), ._C(IC107_7_TO_IC121_4), ._D(IC107_4_TO_IC121_5), ._QA(), ._QB(), ._QC(), ._QD(AZ));

	/* IC122 - LS95 */
	ls95 IC122(._CLK1(SFT_AL), ._CLK2(SFT_AL), ._SER(), ._MODE(LD_SFT_AL), ._A(IC108_12_TO_IC122_2), ._B(IC108_9_TO_IC122_3), ._C(IC108_7_TO_IC122_4), ._D(IC108_4_TO_IC122_5), ._QA(), ._QB(), ._QC(), ._QD(AR));

	/* IC123 - LS95 */
	ls95 IC123(._CLK1(SFT_AL), ._CLK2(SFT_AL), ._SER(), ._MODE(LD_SFT_AL), ._A(IC109_12_TO_IC123_2), ._B(IC109_9_TO_IC123_3), ._C(IC109_7_TO_IC123_4), ._D(IC109_4_TO_IC123_5), ._QA(), ._QB(), ._QC(), ._QD(AG));

	/* IC124 - LS95 */
	ls95 IC124(._CLK1(SFT_AL), ._CLK2(SFT_AL), ._SER(), ._MODE(LD_SFT_AL), ._A(IC110_12_TO_IC124_2), ._B(IC110_9_TO_IC124_3), ._C(IC110_7_TO_IC124_4), ._D(IC110_4_TO_IC124_5), ._QA(), ._QB(), ._QC(), ._QD(AB));

	/* IC136 - LS32 */
	ls32 IC136(._1A(ABHF_AL), ._1B(IC138_8_TO_IC136_2_AND_IC136_5_AND_IC136_10), ._1Y(IC136_3_TO_IC137_13), ._2A(ARHF_AL), ._2B(IC138_8_TO_IC136_2_AND_IC136_5_AND_IC136_10), ._2Y(IC136_6_TO_IC137_5), ._3A(AGHF_AL), ._3B(IC138_8_TO_IC136_2_AND_IC136_5_AND_IC136_10), ._3Y(IC136_8_TO_IC137_9), ._4A(1'b1), ._4B(1'b1), ._4Y());

	/* IC137 - LS10 */
	ls10 IC137(._1A(AB), ._1B(IC139_11_TO_IC137_2_AND_IC137_3_AND_IC137_11), ._1C(IC136_3_TO_IC137_13), ._1Y(AVB), ._2A(IC139_11_TO_IC137_2_AND_IC137_3_AND_IC137_11), ._2B(AR), ._2C(IC136_6_TO_IC137_5), ._2Y(AVR), ._3A(IC136_8_TO_IC137_9), ._3B(AG), ._3C(IC139_11_TO_IC137_2_AND_IC137_3_AND_IC137_11), ._3Y(AVG));

	/* IC138 - LS32 */
	ls32 IC138(._1A(AB), ._1B(AG), ._1Y(IC138_3_TO_IC138_4), ._2A(IC138_3_TO_IC138_4), ._2B(IC138_11_TO_IC138_5), ._2Y(AY_AL), ._3A(KOS1), ._3B(AZ), ._3Y(IC138_8_TO_IC136_2_AND_IC136_5_AND_IC136_10), ._4A(AR), ._4B(AZ), ._4Y(IC138_11_TO_IC138_5));


	/* -> External Shared Logic
	// IC117 - LS04
	// ls04 IC117(._1A(CN1[35]), ._1Y(IC117_2_TO_IC131_1), ._2A(CN1[37]), ._2Y(IC117_3_TO_IC133_4), ._3A(CN1[39]), ._3Y(IC117_6_TO_IC133_9), ._4A(CN1[34]), ._4Y(IC117_8_TO_IC131_11), ._5A(SEL_I_II_AL_A), ._5Y(IC117_10_TO_IC107_1_AND_IC108_1_AND_IC109_1_AND_IC110_1), ._6A(SEL_I_II_AL_B), ._6Y(IC117_12_TO_IC111_1_AND_IC112_1_AND_IC113_1_AND_IC114_1));
	//
	// IC139 - LS00
	// ls00 IC139(._1A(PRIB_AL), ._1B(AY_AL), ._1Y(IC139_3_TO_IC141_2_AND_IC141_3_AND_IC141_11), ._2A(ENB), ._2B(AV6_TICK_AL), ._2Y(IC139_6_TO_IC111_15_AND_IC112_15_AND_IC113_15_AND_IC114_15), ._3A(ENA), ._3B(AV6_TICK_AL), ._3Y(IC139_8_TO_IC107_15_AND_IC108_15_AND_IC109_15_AND_IC110_15), ._4A(BY_AL), ._4B(PRIA_AL), ._4Y(IC139_11_TO_IC137_2_AND_IC137_3_AND_IC137_11));
	*/

endmodule
