/*#########################################################################
#File Name:     ls393_tb.sv
#Description:   SN74LS393N - Dual 4-Bit Decade and Binary Counters test bench.
#    			                      
#Date:          
#Programmer:    Jonathon McEllin, S00150412
#Version:       Rev. 1.00
#
#Notes:         
##########################################################################*/

`timescale 1ps / 1ps
module ls393_tb; 
/*-------------------------- Inputs and Outputs --------------------------*/
	reg    _1A, _1CLR, _2A, _2CLR;
 	wire   _1QA, _1QB, _1QC, _1QD, _2QA, _2QB, _2QC, _2QD;
	
/*--------------------- Instantiate Device Under Test --------------------*/
	ls393 DUT( 
		._1A(_1A),
		._1QA(_1QA),
		._1QB(_1QB),
		._1QC(_1QC),
		._1QD(_1QD),
		._1CLR(_1CLR),
		._2A(_2A),
		._2QA(_2QA),		
		._2QB(_2QB),
		._2QC(_2QC),
		._2QD(_2QD),
		._2CLR(_2CLR)
	);		

/*--------------------------------- Test ---------------------------------*/
	initial begin
		// Reset flip flops
		_1A = 1'b0; _1CLR = 1'b1; _2A = 1'b0; _2CLR = 1'b1;

		// Count up
		#10 _1A = 1'b1;  _1CLR = 1'b0; _2A = 1'b1; _2CLR = 1'b0;
		#10 _1A = 1'b0;  _2A = 1'b0; // 1
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 2
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 3
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 4
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 5
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 6
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 7
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 8
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 9
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 10
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 11
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 12
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 13
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 14
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 15
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 0
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 1
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 2
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 3
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 4
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 5
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 6
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 7
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 8
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 9
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 10
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 11
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 12
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 13
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 14
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 15
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 0
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 1
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 2
		#10 _1A = 1'b1;  _2A = 1'b1;

		// Clear
		#10 _1CLR = 1'b1; _2CLR = 1'b1; // 0
		#10 _1CLR = 1'b0; _2CLR = 1'b0;
		#10 _1A = 1'b0;  _2A = 1'b0; // 1
		#10 _1A = 1'b1;  _2A = 1'b1;
		#10 _1A = 1'b0;  _2A = 1'b0; // 2
		#10 _1A = 1'b1;  _2A = 1'b1;

		#10 $stop;
	end
	
endmodule