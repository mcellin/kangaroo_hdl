/*#########################################################################
#File Name:     ls367_tb.sv
#Description:   M74LS367AP - High-Speed CMOS Logic Hex Buffer/Line Driver,
#    			Three-State Non-Inverting test bench.                        
#
#Date:          
#Programmer:    Jonathon McEllin, S00150412
#Version:       Rev. 1.00
#
#Notes:         
##########################################################################*/

`timescale 1ps / 1ps
module ls367_tb; 
/*-------------------------- Inputs and Outputs --------------------------*/
	reg    _1G, _1A1, _1A2, _1A3, _1A4, _2G, _2A1, _2A2;
 	wire   _1Y1, _1Y2, _1Y3, _1Y4, _2Y1, _2Y2;

/*--------------------- Instantiate Device Under Test --------------------*/
	ls367 DUT( 
		._1G(_1G),
		._1A1(_1A1),
		._1Y1(_1Y1),
		._1A2(_1A2),
		._1Y2(_1Y2),
		._1A3(_1A3),
		._1Y3(_1Y3),
		._1A4(_1A4),		
		._1Y4(_1Y4),
		._2G(_2G),
		._2A1(_2A1),
		._2Y1(_2Y1),		
		._2A2(_2A2),
		._2Y2(_2Y2)
	);

/*--------------------------------- Test ---------------------------------*/
	initial begin
		/*Output Enabled.*/
		_1G = 1'b0; _1A1 = 1'b0; _1A2 = 1'b0; _1A3 = 1'b0; _1A4 = 1'b0; _2G = 1'b0; _2A1 = 1'b0; _2A2 = 1'b0;
		#0 $display("_1G = %b, _1A1 = %b, _1A2 = %b, _1A3 = %b, _1A4 = %b, _2G = %b, _2A1 = %b, _2A2 = %b", _1G, _1A1, _1A2, _1A3, _1A4, _2G, _2A1, _2A2);
		#0 $display("_1Y1 = %b, _1Y2 = %b, _1Y3 = %b, _1Y4 = %b, _2Y1 = %b, _2Y2 = %b", _1Y1, _1Y2, _1Y3, _1Y4, _2Y1, _2Y2);
		
		#10 _1A1 = 1'b1;
		#0 $display("_1G = %b, _1A1 = %b, _1A2 = %b, _1A3 = %b, _1A4 = %b, _2G = %b, _2A1 = %b, _2A2 = %b", _1G, _1A1, _1A2, _1A3, _1A4, _2G, _2A1, _2A2);
		#0 $display("_1Y1 = %b, _1Y2 = %b, _1Y3 = %b, _1Y4 = %b, _2Y1 = %b, _2Y2 = %b", _1Y1, _1Y2, _1Y3, _1Y4, _2Y1, _2Y2);
		
		#10 _1A1 = 1'b0; _1A2 = 1'b1;
		#0 $display("_1G = %b, _1A1 = %b, _1A2 = %b, _1A3 = %b, _1A4 = %b, _2G = %b, _2A1 = %b, _2A2 = %b", _1G, _1A1, _1A2, _1A3, _1A4, _2G, _2A1, _2A2);
		#0 $display("_1Y1 = %b, _1Y2 = %b, _1Y3 = %b, _1Y4 = %b, _2Y1 = %b, _2Y2 = %b", _1Y1, _1Y2, _1Y3, _1Y4, _2Y1, _2Y2);

		#10 _1A2 = 1'b0; _1A3 = 1'b1;
		#0 $display("_1G = %b, _1A1 = %b, _1A2 = %b, _1A3 = %b, _1A4 = %b, _2G = %b, _2A1 = %b, _2A2 = %b", _1G, _1A1, _1A2, _1A3, _1A4, _2G, _2A1, _2A2);
		#0 $display("_1Y1 = %b, _1Y2 = %b, _1Y3 = %b, _1Y4 = %b, _2Y1 = %b, _2Y2 = %b", _1Y1, _1Y2, _1Y3, _1Y4, _2Y1, _2Y2);

		#10 _1A3 = 1'b0; _1A4 = 1'b1;
		#0 $display("_1G = %b, _1A1 = %b, _1A2 = %b, _1A3 = %b, _1A4 = %b, _2G = %b, _2A1 = %b, _2A2 = %b", _1G, _1A1, _1A2, _1A3, _1A4, _2G, _2A1, _2A2);
		#0 $display("_1Y1 = %b, _1Y2 = %b, _1Y3 = %b, _1Y4 = %b, _2Y1 = %b, _2Y2 = %b", _1Y1, _1Y2, _1Y3, _1Y4, _2Y1, _2Y2);

		#10 _1A4 = 1'b0; _2A1 = 1'b1;
		#0 $display("_1G = %b, _1A1 = %b, _1A2 = %b, _1A3 = %b, _1A4 = %b, _2G = %b, _2A1 = %b, _2A2 = %b", _1G, _1A1, _1A2, _1A3, _1A4, _2G, _2A1, _2A2);
		#0 $display("_1Y1 = %b, _1Y2 = %b, _1Y3 = %b, _1Y4 = %b, _2Y1 = %b, _2Y2 = %b", _1Y1, _1Y2, _1Y3, _1Y4, _2Y1, _2Y2);
		
		#10 _2A1 = 1'b0; _2A2 = 1'b1;
		#0 $display("_1G = %b, _1A1 = %b, _1A2 = %b, _1A3 = %b, _1A4 = %b, _2G = %b, _2A1 = %b, _2A2 = %b", _1G, _1A1, _1A2, _1A3, _1A4, _2G, _2A1, _2A2);
		#0 $display("_1Y1 = %b, _1Y2 = %b, _1Y3 = %b, _1Y4 = %b, _2Y1 = %b, _2Y2 = %b", _1Y1, _1Y2, _1Y3, _1Y4, _2Y1, _2Y2);

		/*Output Disabled. Check for high impedence*/
		#10 _1G = 1'b1; _2G = 1'b1; _2A2 = 1'b0;
		#0 $display("_1G = %b, _1A1 = %b, _1A2 = %b, _1A3 = %b, _1A4 = %b, _2G = %b, _2A1 = %b, _2A2 = %b", _1G, _1A1, _1A2, _1A3, _1A4, _2G, _2A1, _2A2);
		#0 $display("_1Y1 = %b, _1Y2 = %b, _1Y3 = %b, _1Y4 = %b, _2Y1 = %b, _2Y2 = %b", _1Y1, _1Y2, _1Y3, _1Y4, _2Y1, _2Y2);
		
		#10 _1A1 = 1'b1;
		#0 $display("_1G = %b, _1A1 = %b, _1A2 = %b, _1A3 = %b, _1A4 = %b, _2G = %b, _2A1 = %b, _2A2 = %b", _1G, _1A1, _1A2, _1A3, _1A4, _2G, _2A1, _2A2);
		#0 $display("_1Y1 = %b, _1Y2 = %b, _1Y3 = %b, _1Y4 = %b, _2Y1 = %b, _2Y2 = %b", _1Y1, _1Y2, _1Y3, _1Y4, _2Y1, _2Y2);
		
		#10 _1A1 = 1'b0; _1A2 = 1'b1;
		#0 $display("_1G = %b, _1A1 = %b, _1A2 = %b, _1A3 = %b, _1A4 = %b, _2G = %b, _2A1 = %b, _2A2 = %b", _1G, _1A1, _1A2, _1A3, _1A4, _2G, _2A1, _2A2);
		#0 $display("_1Y1 = %b, _1Y2 = %b, _1Y3 = %b, _1Y4 = %b, _2Y1 = %b, _2Y2 = %b", _1Y1, _1Y2, _1Y3, _1Y4, _2Y1, _2Y2);

		#10 _1A2 = 1'b0; _1A3 = 1'b1;
		#0 $display("_1G = %b, _1A1 = %b, _1A2 = %b, _1A3 = %b, _1A4 = %b, _2G = %b, _2A1 = %b, _2A2 = %b", _1G, _1A1, _1A2, _1A3, _1A4, _2G, _2A1, _2A2);
		#0 $display("_1Y1 = %b, _1Y2 = %b, _1Y3 = %b, _1Y4 = %b, _2Y1 = %b, _2Y2 = %b", _1Y1, _1Y2, _1Y3, _1Y4, _2Y1, _2Y2);

		#10 _1A3 = 1'b0; _1A4 = 1'b1;
		#0 $display("_1G = %b, _1A1 = %b, _1A2 = %b, _1A3 = %b, _1A4 = %b, _2G = %b, _2A1 = %b, _2A2 = %b", _1G, _1A1, _1A2, _1A3, _1A4, _2G, _2A1, _2A2);
		#0 $display("_1Y1 = %b, _1Y2 = %b, _1Y3 = %b, _1Y4 = %b, _2Y1 = %b, _2Y2 = %b", _1Y1, _1Y2, _1Y3, _1Y4, _2Y1, _2Y2);

		#10 _1A4 = 1'b0; _2A1 = 1'b1;
		#0 $display("_1G = %b, _1A1 = %b, _1A2 = %b, _1A3 = %b, _1A4 = %b, _2G = %b, _2A1 = %b, _2A2 = %b", _1G, _1A1, _1A2, _1A3, _1A4, _2G, _2A1, _2A2);
		#0 $display("_1Y1 = %b, _1Y2 = %b, _1Y3 = %b, _1Y4 = %b, _2Y1 = %b, _2Y2 = %b", _1Y1, _1Y2, _1Y3, _1Y4, _2Y1, _2Y2);
		
		#10 _2A1 = 1'b0; _2A2 = 1'b1;
		#0 $display("_1G = %b, _1A1 = %b, _1A2 = %b, _1A3 = %b, _1A4 = %b, _2G = %b, _2A1 = %b, _2A2 = %b", _1G, _1A1, _1A2, _1A3, _1A4, _2G, _2A1, _2A2);
		#0 $display("_1Y1 = %b, _1Y2 = %b, _1Y3 = %b, _1Y4 = %b, _2Y1 = %b, _2Y2 = %b", _1Y1, _1Y2, _1Y3, _1Y4, _2Y1, _2Y2);

		#10 $stop;
	end
	
endmodule